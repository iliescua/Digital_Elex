#Creating an NMOS inverter
.model nmod NMOS KP=346U VTO=1.18V

VDD 1 0 DC 5V
R1 1 2 100K
VA 3 0 DC 5V
M1 2 3 0 0 nmod W=4U L=2U

.dc VA 0 5 0.01
