#Creating the TTL inverter for the prelab and getting its measurements
.model npnt NPN BF=100 IS=1.8f
.model diode D IS=1pA n=1.8 BV=75

VCC 1 0 DC 5V
RC 1 2 3.9k
RB 1 3 3.9k
VA 4 0 5V
Q1 5 3 4 npnt
Q2 2 5 0 npnt


.dc VA 0 5 0.001
.end
